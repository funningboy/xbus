

`define DEF_C_RW_WIDTH    1
`define DEF_C_REQ_WIDTH   1
`define DEF_C_ACK_WIDTH   1
`define DEF_C_ADDR_WIDTH  14
`define DEF_C_BE_WIDTH    4
`define DEF_C_RDATA_WIDTH 32
`define DEF_C_WDATA_WIDTH 32
`define DEF_C_CLK_PERIOD  5
